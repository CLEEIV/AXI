module Interconnect (
    //----- Global -----//
    input  ACLK   ,
    input  ARESETn,
    //----- Master 0 -----//
    // Write adress
    input  [3:0]  m0_axi_awid   ,
    input  [31:0] m0_axi_awaddr ,
    input  [7:0]  m0_axi_awlen  ,
    input  [2:0]  m0_axi_awsize ,
    input  [1:0]  m0_axi_awburst,
    input         m0_axi_awvalid,
    output        m0_axi_awready,
    // Write data
    input  [31:0] m0_axi_wdata  ,
    input  [3:0]  m0_axi_wstrb  ,
    input         m0_axi_wlast  ,
    input         m0_axi_wvalid ,
    output        m0_axi_wready ,
    // Write response
    output [3:0]  m0_axi_bid    ,
    output [1:0]  m0_axi_bresp  ,
    output        m0_axi_bvalid ,
    input         m0_axi_bready ,
    // Read address
    input  [3:0]  m0_axi_arid   ,
    input  [31:0] m0_axi_araddr ,
    input  [7:0]  m0_axi_arlen  ,
    input  [2:0]  m0_axi_arsize ,
    input  [1:0]  m0_axi_arburst,
    input         m0_axi_arvalid,
    output        m0_axi_arready,
    // Read data
    output [3:0]  m0_axi_rid    ,
    output [31:0] m0_axi_rdata  ,
    output [1:0]  m0_axi_rresp  ,
    output        m0_axi_rlast  ,
    output        m0_axi_rvalid ,
    input         m0_axi_rready ,
    //----- Master 1 -----//
    // Write adress
    input  [3:0]  m1_axi_awid   ,
    input  [31:0] m1_axi_awaddr ,
    input  [7:0]  m1_axi_awlen  ,
    input  [2:0]  m1_axi_awsize ,
    input  [1:0]  m1_axi_awburst,
    input         m1_axi_awvalid,
    output        m1_axi_awready,
    // Write data
    input  [31:0] m1_axi_wdata  ,
    input  [3:0]  m1_axi_wstrb  ,
    input         m1_axi_wlast  ,
    input         m1_axi_wvalid ,
    output        m1_axi_wready ,
    // Write response
    output [3:0]  m1_axi_bid    ,
    output [1:0]  m1_axi_bresp  ,
    output        m1_axi_bvalid ,
    input         m1_axi_bready ,
    // Read address
    input  [3:0]  m1_axi_arid   ,
    input  [31:0] m1_axi_araddr ,
    input  [7:0]  m1_axi_arlen  ,
    input  [2:0]  m1_axi_arsize ,
    input  [1:0]  m1_axi_arburst,
    input         m1_axi_arvalid,
    output        m1_axi_arready,
    // Read data
    output [3:0]  m1_axi_rid    ,
    output [31:0] m1_axi_rdata  ,
    output [1:0]  m1_axi_rresp  ,
    output        m1_axi_rlast  ,
    output        m1_axi_rvalid ,
    input         m1_axi_rready ,
    //----- Master 2 -----//
    // Write adress
    input  [3:0]  m2_axi_awid   ,
    input  [31:0] m2_axi_awaddr ,
    input  [7:0]  m2_axi_awlen  ,
    input  [2:0]  m2_axi_awsize ,
    input  [1:0]  m2_axi_awburst,
    input         m2_axi_awvalid,
    output        m2_axi_awready,
    // Write data
    input  [31:0] m2_axi_wdata  ,
    input  [3:0]  m2_axi_wstrb  ,
    input         m2_axi_wlast  ,
    input         m2_axi_wvalid ,
    output        m2_axi_wready ,
    // Write response
    output [3:0]  m2_axi_bid    ,
    output [1:0]  m2_axi_bresp  ,
    output        m2_axi_bvalid ,
    input         m2_axi_bready ,
    // Read address
    input  [3:0]  m2_axi_arid   ,
    input  [31:0] m2_axi_araddr ,
    input  [7:0]  m2_axi_arlen  ,
    input  [2:0]  m2_axi_arsize ,
    input  [1:0]  m2_axi_arburst,
    input         m2_axi_arvalid,
    output        m2_axi_arready,
    // Read data
    output [3:0]  m2_axi_rid    ,
    output [31:0] m2_axi_rdata  ,
    output [1:0]  m2_axi_rresp  ,
    output        m2_axi_rlast  ,
    output        m2_axi_rvalid ,
    input         m2_axi_rready ,
    //----- Master 3 -----//
    // Write adress
    input  [3:0]  m3_axi_awid   ,
    input  [31:0] m3_axi_awaddr ,
    input  [7:0]  m3_axi_awlen  ,
    input  [2:0]  m3_axi_awsize ,
    input  [1:0]  m3_axi_awburst,
    input         m3_axi_awvalid,
    output        m3_axi_awready,
    // Write data
    input  [31:0] m3_axi_wdata  ,
    input  [3:0]  m3_axi_wstrb  ,
    input         m3_axi_wlast  ,
    input         m3_axi_wvalid ,
    output        m3_axi_wready ,
    // Write response
    output [3:0]  m3_axi_bid    ,
    output [1:0]  m3_axi_bresp  ,
    output        m3_axi_bvalid ,
    input         m3_axi_bready ,
    // Read address
    input  [3:0]  m3_axi_arid   ,
    input  [31:0] m3_axi_araddr ,
    input  [7:0]  m3_axi_arlen  ,
    input  [2:0]  m3_axi_arsize ,
    input  [1:0]  m3_axi_arburst,
    input         m3_axi_arvalid,
    output        m3_axi_arready,
    // Read data
    output [3:0]  m3_axi_rid    ,
    output [31:0] m3_axi_rdata  ,
    output [1:0]  m3_axi_rresp  ,
    output        m3_axi_rlast  ,
    output        m3_axi_rvalid ,
    input         m3_axi_rready ,
    //----- Slave 0 -----//
    // Write adress
    output [3:0]  s0_axi_awid   ,
    output [31:0] s0_axi_awaddr ,
    output [7:0]  s0_axi_awlen  ,
    output [2:0]  s0_axi_awsize ,
    output [1:0]  s0_axi_awburst,
    output        s0_axi_awvalid,
    input         s0_axi_awready,
    // Write data
    output [31:0] s0_axi_wdata  ,
    output [3:0]  s0_axi_wstrb  ,
    output        s0_axi_wlast  ,
    output        s0_axi_wvalid ,
    input         s0_axi_wready ,
    // Write response
    input  [3:0]  s0_axi_bid    ,
    input  [1:0]  s0_axi_bresp  ,
    input         s0_axi_bvalid ,
    output        s0_axi_bready ,
    // Read address
    output [3:0]  s0_axi_arid   ,
    output [31:0] s0_axi_araddr ,
    output [7:0]  s0_axi_arlen  ,
    output [2:0]  s0_axi_arsize ,
    output [1:0]  s0_axi_arburst,
    output        s0_axi_arvalid,
    input         s0_axi_arready,
    // Read data
    input  [3:0]  s0_axi_rid    ,
    input  [31:0] s0_axi_rdata  ,
    input  [1:0]  s0_axi_rresp  ,
    input         s0_axi_rlast  ,
    input         s0_axi_rvalid ,
    output        s0_axi_rready ,
    //----- Slave 1 -----//
    // Write adress
    output [3:0]  s1_axi_awid   ,
    output [31:0] s1_axi_awaddr ,
    output [7:0]  s1_axi_awlen  ,
    output [2:0]  s1_axi_awsize ,
    output [1:0]  s1_axi_awburst,
    output        s1_axi_awvalid,
    input         s1_axi_awready,
    // Write data
    output [31:0] s1_axi_wdata  ,
    output [3:0]  s1_axi_wstrb  ,
    output        s1_axi_wlast  ,
    output        s1_axi_wvalid ,
    input         s1_axi_wready ,
    // Write response
    input  [3:0]  s1_axi_bid    ,
    input  [1:0]  s1_axi_bresp  ,
    input         s1_axi_bvalid ,
    output        s1_axi_bready ,
    // Read address
    output [3:0]  s1_axi_arid   ,
    output [31:0] s1_axi_araddr ,
    output [7:0]  s1_axi_arlen  ,
    output [2:0]  s1_axi_arsize ,
    output [1:0]  s1_axi_arburst,
    output        s1_axi_arvalid,
    input         s1_axi_arready,
    // Read data
    input  [3:0]  s1_axi_rid    ,
    input  [31:0] s1_axi_rdata  ,
    input  [1:0]  s1_axi_rresp  ,
    input         s1_axi_rlast  ,
    input         s1_axi_rvalid ,
    output        s1_axi_rready ,
    //----- Slave 2 -----//
    // Write adress
    output [3:0]  s2_axi_awid   ,
    output [31:0] s2_axi_awaddr ,
    output [7:0]  s2_axi_awlen  ,
    output [2:0]  s2_axi_awsize ,
    output [1:0]  s2_axi_awburst,
    output        s2_axi_awvalid,
    input         s2_axi_awready,
    // Write data
    output [31:0] s2_axi_wdata  ,
    output [3:0]  s2_axi_wstrb  ,
    output        s2_axi_wlast  ,
    output        s2_axi_wvalid ,
    input         s2_axi_wready ,
    // Write response
    input  [3:0]  s2_axi_bid    ,
    input  [1:0]  s2_axi_bresp  ,
    input         s2_axi_bvalid ,
    output        s2_axi_bready ,
    // Read address
    output [3:0]  s2_axi_arid   ,
    output [31:0] s2_axi_araddr ,
    output [7:0]  s2_axi_arlen  ,
    output [2:0]  s2_axi_arsize ,
    output [1:0]  s2_axi_arburst,
    output        s2_axi_arvalid,
    input         s2_axi_arready,
    // Read data
    input  [3:0]  s2_axi_rid    ,
    input  [31:0] s2_axi_rdata  ,
    input  [1:0]  s2_axi_rresp  ,
    input         s2_axi_rlast  ,
    input         s2_axi_rvalid ,
    output        s2_axi_rready ,
    //----- Slave 3 -----//
    // Write adress
    output [3:0]  s3_axi_awid   ,
    output [31:0] s3_axi_awaddr ,
    output [7:0]  s3_axi_awlen  ,
    output [2:0]  s3_axi_awsize ,
    output [1:0]  s3_axi_awburst,
    output        s3_axi_awvalid,
    input         s3_axi_awready,
    // Write data
    output [31:0] s3_axi_wdata  ,
    output [3:0]  s3_axi_wstrb  ,
    output        s3_axi_wlast  ,
    output        s3_axi_wvalid ,
    input         s3_axi_wready ,
    // Write response
    input  [3:0]  s3_axi_bid    ,
    input  [1:0]  s3_axi_bresp  ,
    input         s3_axi_bvalid ,
    output        s3_axi_bready ,
    // Read address
    output [3:0]  s3_axi_arid   ,
    output [31:0] s3_axi_araddr ,
    output [7:0]  s3_axi_arlen  ,
    output [2:0]  s3_axi_arsize ,
    output [1:0]  s3_axi_arburst,
    output        s3_axi_arvalid,
    input         s3_axi_arready,
    // Read data
    input  [3:0]  s3_axi_rid    ,
    input  [31:0] s3_axi_rdata  ,
    input  [1:0]  s3_axi_rresp  ,
    input         s3_axi_rlast  ,
    input         s3_axi_rvalid ,
    output        s3_axi_rready 
);
wire m0_read_accept ;
wire m1_read_accept ;
wire m2_read_accept ;
wire m3_read_accept ;
wire m0_write_accept;
wire m1_write_accept;
wire m2_write_accept;
wire m3_write_accept;
//----- Master_MUX to Slave_MUX -----//
// Write address
wire        m_awready;
wire [3:0]  s_awid   ;
wire [31:0] s_awaddr ;
wire [7:0]  s_awlen  ;
wire [2:0]  s_awsize ;
wire [1:0]  s_awburst;
wire        s_awvalid;
// Write data
wire        m_wready ;
wire [31:0] s_wdata  ;
wire [3:0]  s_wstrb  ;
wire        s_wlast  ;
wire        s_wvalid ;
// Write response
wire [3:0]  m_bid    ;
wire [1:0]  m_bresp  ;
wire        m_bvalid ;
wire        s_bready ;
// Read address
wire        m_arready;
wire [3:0]  s_arid   ;
wire [31:0] s_araddr ;
wire [7:0]  s_arlen  ;
wire [2:0]  s_arsize ;
wire [1:0]  s_arburst;
wire        s_arvalid;
// Read data
wire [3:0]  m_rid    ;
wire [31:0] m_rdata  ;
wire [1:0]  m_rresp  ;
wire        m_rlast  ;
wire        m_rvalid ;
wire        s_rready ;
Arbiter_R Arbiter_R (
    .aclk           ( ACLK           ),
    .aresetn        ( ARESETn        ),
    .m0_arvalid     ( m0_axi_arvalid ),
    .m0_rready      ( m0_axi_rready  ),
    .m1_arvalid     ( m1_axi_arvalid ),
    .m1_rready      ( m1_axi_rready  ),
    .m2_arvalid     ( m2_axi_arvalid ),
    .m2_rready      ( m2_axi_rready  ),
    .m3_arvalid     ( m3_axi_arvalid ),
    .m3_rready      ( m3_axi_rready  ),
    .m_rvalid       ( m_rvalid       ),
    .m_rlast        ( m_rlast        ),
    .m0_read_accept ( m0_read_accept ),
    .m1_read_accept ( m1_read_accept ),
    .m2_read_accept ( m2_read_accept ),
    .m3_read_accept ( m3_read_accept ) 
);
Arbiter_W Arbiter_W (
    .aclk            ( ACLK            ),
    .aresetn         ( ARESETn         ),
    .m0_awvalid      ( m0_axi_awvalid  ),
    .m0_wvalid       ( m0_axi_wvalid   ),
    .m0_bready       ( m0_axi_bready   ),
    .m1_awvalid      ( m1_axi_awvalid  ),
    .m1_wvalid       ( m1_axi_wvalid   ),
    .m1_bready       ( m1_axi_bready   ),
    .m2_awvalid      ( m2_axi_awvalid  ),
    .m2_wvalid       ( m2_axi_wvalid   ),
    .m2_bready       ( m2_axi_bready   ),
    .m3_awvalid      ( m3_axi_awvalid  ),
    .m3_wvalid       ( m3_axi_wvalid   ),
    .m3_bready       ( m3_axi_bready   ),
    .m_awready       ( m_awready       ),
    .m_wready        ( m_wready        ),
    .m_bvalid        ( m_bvalid        ),
    .m0_write_accept ( m0_write_accept ),
    .m1_write_accept ( m1_write_accept ),
    .m2_write_accept ( m2_write_accept ),
    .m3_write_accept ( m3_write_accept ) 
);
Master_Mux_R Master_Mux_R (
    .aclk           ( ACLK            ),
    .aresetn        ( ARESETn         ),
    .m0_axi_arid    ( m0_axi_arid     ),
    .m0_axi_araddr  ( m0_axi_araddr   ),
    .m0_axi_arlen   ( m0_axi_arlen    ),
    .m0_axi_arsize  ( m0_axi_arsize   ),
    .m0_axi_arburst ( m0_axi_arburst  ),
    .m0_axi_arvalid ( m0_axi_arvalid  ),
    .m0_axi_arready ( m0_axi_arready  ),
    .m0_axi_rid     ( m0_axi_rid      ),
    .m0_axi_rdata   ( m0_axi_rdata    ),
    .m0_axi_rresp   ( m0_axi_rresp    ),
    .m0_axi_rlast   ( m0_axi_rlast    ),
    .m0_axi_rvalid  ( m0_axi_rvalid   ),
    .m0_axi_rready  ( m0_axi_rready   ),
    .m1_axi_arid    ( m1_axi_arid     ),
    .m1_axi_araddr  ( m1_axi_araddr   ),
    .m1_axi_arlen   ( m1_axi_arlen    ),
    .m1_axi_arsize  ( m1_axi_arsize   ),
    .m1_axi_arburst ( m1_axi_arburst  ),
    .m1_axi_arvalid ( m1_axi_arvalid  ),
    .m1_axi_arready ( m1_axi_arready  ),
    .m1_axi_rid     ( m1_axi_rid      ),
    .m1_axi_rdata   ( m1_axi_rdata    ),
    .m1_axi_rresp   ( m1_axi_rresp    ),
    .m1_axi_rlast   ( m1_axi_rlast    ),
    .m1_axi_rvalid  ( m1_axi_rvalid   ),
    .m1_axi_rready  ( m1_axi_rready   ),
    .m2_axi_arid    ( m2_axi_arid     ),
    .m2_axi_araddr  ( m2_axi_araddr   ),
    .m2_axi_arlen   ( m2_axi_arlen    ),
    .m2_axi_arsize  ( m2_axi_arsize   ),
    .m2_axi_arburst ( m2_axi_arburst  ),
    .m2_axi_arvalid ( m2_axi_arvalid  ),
    .m2_axi_arready ( m2_axi_arready  ),
    .m2_axi_rid     ( m2_axi_rid      ),
    .m2_axi_rdata   ( m2_axi_rdata    ),
    .m2_axi_rresp   ( m2_axi_rresp    ),
    .m2_axi_rlast   ( m2_axi_rlast    ),
    .m2_axi_rvalid  ( m2_axi_rvalid   ),
    .m2_axi_rready  ( m2_axi_rready   ),
    .m3_axi_arid    ( m3_axi_arid     ),
    .m3_axi_araddr  ( m3_axi_araddr   ),
    .m3_axi_arlen   ( m3_axi_arlen    ),
    .m3_axi_arsize  ( m3_axi_arsize   ),
    .m3_axi_arburst ( m3_axi_arburst  ),
    .m3_axi_arvalid ( m3_axi_arvalid  ),
    .m3_axi_arready ( m3_axi_arready  ),
    .m3_axi_rid     ( m3_axi_rid      ),
    .m3_axi_rdata   ( m3_axi_rdata    ),
    .m3_axi_rresp   ( m3_axi_rresp    ),
    .m3_axi_rlast   ( m3_axi_rlast    ),
    .m3_axi_rvalid  ( m3_axi_rvalid   ),
    .m3_axi_rready  ( m3_axi_rready   ),
    .s_arid         ( s_arid          ),
    .s_araddr       ( s_araddr        ),
    .s_arlen        ( s_arlen         ),
    .s_arsize       ( s_arsize        ),
    .s_arburst      ( s_arburst       ),
    .s_arvalid      ( s_arvalid       ),
    .s_rready       ( s_rready        ),
    .m_arready      ( m_arready       ),
    .m_rid          ( m_rid           ),
    .m_rdata        ( m_rdata         ),
    .m_rresp        ( m_rresp         ),
    .m_rlast        ( m_rlast         ),
    .m_rvalid       ( m_rvalid        ),
    .m0_read_accept ( m0_read_accept  ),
    .m1_read_accept ( m1_read_accept  ),
    .m2_read_accept ( m2_read_accept  ),
    .m3_read_accept ( m3_read_accept  )
);
Master_Mux_W Master_Mux_W (
    .aclk            ( ACLK            ),
    .aresetn         ( ARESETn         ),
    .m0_axi_awid     ( m0_axi_awid     ),
    .m0_axi_awaddr   ( m0_axi_awaddr   ),
    .m0_axi_awlen    ( m0_axi_awlen    ),
    .m0_axi_awsize   ( m0_axi_awsize   ),
    .m0_axi_awburst  ( m0_axi_awburst  ),
    .m0_axi_awvalid  ( m0_axi_awvalid  ),
    .m0_axi_awready  ( m0_axi_awready  ),
    .m0_axi_wdata    ( m0_axi_wdata    ),
    .m0_axi_wstrb    ( m0_axi_wstrb    ),
    .m0_axi_wlast    ( m0_axi_wlast    ),
    .m0_axi_wvalid   ( m0_axi_wvalid   ),
    .m0_axi_wready   ( m0_axi_wready   ),
    .m0_axi_bid      ( m0_axi_bid      ),
    .m0_axi_bresp    ( m0_axi_bresp    ),
    .m0_axi_bvalid   ( m0_axi_bvalid   ),
    .m0_axi_bready   ( m0_axi_bready   ),
    .m1_axi_awid     ( m1_axi_awid     ),
    .m1_axi_awaddr   ( m1_axi_awaddr   ),
    .m1_axi_awlen    ( m1_axi_awlen    ),
    .m1_axi_awsize   ( m1_axi_awsize   ),
    .m1_axi_awburst  ( m1_axi_awburst  ),
    .m1_axi_awvalid  ( m1_axi_awvalid  ),
    .m1_axi_awready  ( m1_axi_awready  ),
    .m1_axi_wdata    ( m1_axi_wdata    ),
    .m1_axi_wstrb    ( m1_axi_wstrb    ),
    .m1_axi_wlast    ( m1_axi_wlast    ),
    .m1_axi_wvalid   ( m1_axi_wvalid   ),
    .m1_axi_wready   ( m1_axi_wready   ),
    .m1_axi_bid      ( m1_axi_bid      ),
    .m1_axi_bresp    ( m1_axi_bresp    ),
    .m1_axi_bvalid   ( m1_axi_bvalid   ),
    .m1_axi_bready   ( m1_axi_bready   ),
    .m2_axi_awid     ( m2_axi_awid     ),
    .m2_axi_awaddr   ( m2_axi_awaddr   ),
    .m2_axi_awlen    ( m2_axi_awlen    ),
    .m2_axi_awsize   ( m2_axi_awsize   ),
    .m2_axi_awburst  ( m2_axi_awburst  ),
    .m2_axi_awvalid  ( m2_axi_awvalid  ),
    .m2_axi_awready  ( m2_axi_awready  ),
    .m2_axi_wdata    ( m2_axi_wdata    ),
    .m2_axi_wstrb    ( m2_axi_wstrb    ),
    .m2_axi_wlast    ( m2_axi_wlast    ),
    .m2_axi_wvalid   ( m2_axi_wvalid   ),
    .m2_axi_wready   ( m2_axi_wready   ),
    .m2_axi_bid      ( m2_axi_bid      ),
    .m2_axi_bresp    ( m2_axi_bresp    ),
    .m2_axi_bvalid   ( m2_axi_bvalid   ),
    .m2_axi_bready   ( m2_axi_bready   ),
    .m3_axi_awid     ( m3_axi_awid     ),
    .m3_axi_awaddr   ( m3_axi_awaddr   ),
    .m3_axi_awlen    ( m3_axi_awlen    ),
    .m3_axi_awsize   ( m3_axi_awsize   ),
    .m3_axi_awburst  ( m3_axi_awburst  ),
    .m3_axi_awvalid  ( m3_axi_awvalid  ),
    .m3_axi_awready  ( m3_axi_awready  ),
    .m3_axi_wdata    ( m3_axi_wdata    ),
    .m3_axi_wstrb    ( m3_axi_wstrb    ),
    .m3_axi_wlast    ( m3_axi_wlast    ),
    .m3_axi_wvalid   ( m3_axi_wvalid   ),
    .m3_axi_wready   ( m3_axi_wready   ),
    .m3_axi_bid      ( m3_axi_bid      ),
    .m3_axi_bresp    ( m3_axi_bresp    ),
    .m3_axi_bvalid   ( m3_axi_bvalid   ),
    .m3_axi_bready   ( m3_axi_bready   ),
    .s_awid          ( s_awid          ),
    .s_awaddr        ( s_awaddr        ),
    .s_awlen         ( s_awlen         ),
    .s_awsize        ( s_awsize        ),
    .s_awburst       ( s_awburst       ),
    .s_awvalid       ( s_awvalid       ),
    .s_wdata         ( s_wdata         ),
    .s_wstrb         ( s_wstrb         ),
    .s_wlast         ( s_wlast         ),
    .s_wvalid        ( s_wvalid        ),
    .s_bready        ( s_bready        ),
    .m_awready       ( m_awready       ),
    .m_wready        ( m_wready        ),
    .m_bid           ( m_bid           ),
    .m_bresp         ( m_bresp         ),
    .m_bvalid        ( m_bvalid        ),
    .m0_write_accept ( m0_write_accept ),
    .m1_write_accept ( m1_write_accept ),
    .m2_write_accept ( m2_write_accept ),
    .m3_write_accept ( m3_write_accept )
);
Slave_Mux_R Slave_Mux_R (
    .aclk           ( ACLK           ),
    .aresetn        ( ARESETn        ),
    .s0_axi_arid    ( s0_axi_arid    ),
    .s0_axi_araddr  ( s0_axi_araddr  ),
    .s0_axi_arlen   ( s0_axi_arlen   ),
    .s0_axi_arsize  ( s0_axi_arsize  ),
    .s0_axi_arburst ( s0_axi_arburst ),
    .s0_axi_arvalid ( s0_axi_arvalid ),
    .s0_axi_arready ( s0_axi_arready ),
    .s0_axi_rid     ( s0_axi_rid     ),
    .s0_axi_rdata   ( s0_axi_rdata   ),
    .s0_axi_rresp   ( s0_axi_rresp   ),
    .s0_axi_rlast   ( s0_axi_rlast   ),
    .s0_axi_rvalid  ( s0_axi_rvalid  ),
    .s0_axi_rready  ( s0_axi_rready  ),
    .s1_axi_arid    ( s1_axi_arid    ),
    .s1_axi_araddr  ( s1_axi_araddr  ),
    .s1_axi_arlen   ( s1_axi_arlen   ),
    .s1_axi_arsize  ( s1_axi_arsize  ),
    .s1_axi_arburst ( s1_axi_arburst ),
    .s1_axi_arvalid ( s1_axi_arvalid ),
    .s1_axi_arready ( s1_axi_arready ),
    .s1_axi_rid     ( s1_axi_rid     ),
    .s1_axi_rdata   ( s1_axi_rdata   ),
    .s1_axi_rresp   ( s1_axi_rresp   ),
    .s1_axi_rlast   ( s1_axi_rlast   ),
    .s1_axi_rvalid  ( s1_axi_rvalid  ),
    .s1_axi_rready  ( s1_axi_rready  ),
    .s2_axi_arid    ( s2_axi_arid    ),
    .s2_axi_araddr  ( s2_axi_araddr  ),
    .s2_axi_arlen   ( s2_axi_arlen   ),
    .s2_axi_arsize  ( s2_axi_arsize  ),
    .s2_axi_arburst ( s2_axi_arburst ),
    .s2_axi_arvalid ( s2_axi_arvalid ),
    .s2_axi_arready ( s2_axi_arready ),
    .s2_axi_rid     ( s2_axi_rid     ),
    .s2_axi_rdata   ( s2_axi_rdata   ),
    .s2_axi_rresp   ( s2_axi_rresp   ),
    .s2_axi_rlast   ( s2_axi_rlast   ),
    .s2_axi_rvalid  ( s2_axi_rvalid  ),
    .s2_axi_rready  ( s2_axi_rready  ),
    .s3_axi_arid    ( s3_axi_arid    ),
    .s3_axi_araddr  ( s3_axi_araddr  ),
    .s3_axi_arlen   ( s3_axi_arlen   ),
    .s3_axi_arsize  ( s3_axi_arsize  ),
    .s3_axi_arburst ( s3_axi_arburst ),
    .s3_axi_arvalid ( s3_axi_arvalid ),
    .s3_axi_arready ( s3_axi_arready ),
    .s3_axi_rid     ( s3_axi_rid     ),
    .s3_axi_rdata   ( s3_axi_rdata   ),
    .s3_axi_rresp   ( s3_axi_rresp   ),
    .s3_axi_rlast   ( s3_axi_rlast   ),
    .s3_axi_rvalid  ( s3_axi_rvalid  ),
    .s3_axi_rready  ( s3_axi_rready  ),
    .m_arready      ( m_arready      ),
    .m_rid          ( m_rid          ),
    .m_rdata        ( m_rdata        ),
    .m_rresp        ( m_rresp        ),
    .m_rlast        ( m_rlast        ),
    .m_rvalid       ( m_rvalid       ),
    .s_arid         ( s_arid         ),
    .s_araddr       ( s_araddr       ),
    .s_arlen        ( s_arlen        ),
    .s_arsize       ( s_arsize       ),
    .s_arburst      ( s_arburst      ),
    .s_arvalid      ( s_arvalid      ),
    .s_rready       ( s_rready       )
);
Slave_Mux_W Slave_Mux_W (
    .aclk           ( ACLK           ),
    .aresetn        ( ARESETn        ),
    .s0_axi_awid    ( s0_axi_awid    ),
    .s0_axi_awaddr  ( s0_axi_awaddr  ),
    .s0_axi_awlen   ( s0_axi_awlen   ),
    .s0_axi_awsize  ( s0_axi_awsize  ),
    .s0_axi_awburst ( s0_axi_awburst ),
    .s0_axi_awvalid ( s0_axi_awvalid ),
    .s0_axi_awready ( s0_axi_awready ),
    .s0_axi_wdata   ( s0_axi_wdata   ),
    .s0_axi_wstrb   ( s0_axi_wstrb   ),
    .s0_axi_wlast   ( s0_axi_wlast   ),
    .s0_axi_wvalid  ( s0_axi_wvalid  ),
    .s0_axi_wready  ( s0_axi_wready  ),
    .s0_axi_bid     ( s0_axi_bid     ),
    .s0_axi_bresp   ( s0_axi_bresp   ),
    .s0_axi_bvalid  ( s0_axi_bvalid  ),
    .s0_axi_bready  ( s0_axi_bready  ),
    .s1_axi_awid    ( s1_axi_awid    ),
    .s1_axi_awaddr  ( s1_axi_awaddr  ),
    .s1_axi_awlen   ( s1_axi_awlen   ),
    .s1_axi_awsize  ( s1_axi_awsize  ),
    .s1_axi_awburst ( s1_axi_awburst ),
    .s1_axi_awvalid ( s1_axi_awvalid ),
    .s1_axi_awready ( s1_axi_awready ),
    .s1_axi_wdata   ( s1_axi_wdata   ),
    .s1_axi_wstrb   ( s1_axi_wstrb   ),
    .s1_axi_wlast   ( s1_axi_wlast   ),
    .s1_axi_wvalid  ( s1_axi_wvalid  ),
    .s1_axi_wready  ( s1_axi_wready  ),
    .s1_axi_bid     ( s1_axi_bid     ),
    .s1_axi_bresp   ( s1_axi_bresp   ),
    .s1_axi_bvalid  ( s1_axi_bvalid  ),
    .s1_axi_bready  ( s1_axi_bready  ),
    .s2_axi_awid    ( s2_axi_awid    ),
    .s2_axi_awaddr  ( s2_axi_awaddr  ),
    .s2_axi_awlen   ( s2_axi_awlen   ),
    .s2_axi_awsize  ( s2_axi_awsize  ),
    .s2_axi_awburst ( s2_axi_awburst ),
    .s2_axi_awvalid ( s2_axi_awvalid ),
    .s2_axi_awready ( s2_axi_awready ),
    .s2_axi_wdata   ( s2_axi_wdata   ),
    .s2_axi_wstrb   ( s2_axi_wstrb   ),
    .s2_axi_wlast   ( s2_axi_wlast   ),
    .s2_axi_wvalid  ( s2_axi_wvalid  ),
    .s2_axi_wready  ( s2_axi_wready  ),
    .s2_axi_bid     ( s2_axi_bid     ),
    .s2_axi_bresp   ( s2_axi_bresp   ),
    .s2_axi_bvalid  ( s2_axi_bvalid  ),
    .s2_axi_bready  ( s2_axi_bready  ),
    .s3_axi_awid    ( s3_axi_awid    ),
    .s3_axi_awaddr  ( s3_axi_awaddr  ),
    .s3_axi_awlen   ( s3_axi_awlen   ),
    .s3_axi_awsize  ( s3_axi_awsize  ),
    .s3_axi_awburst ( s3_axi_awburst ),
    .s3_axi_awvalid ( s3_axi_awvalid ),
    .s3_axi_awready ( s3_axi_awready ),
    .s3_axi_wdata   ( s3_axi_wdata   ),
    .s3_axi_wstrb   ( s3_axi_wstrb   ),
    .s3_axi_wlast   ( s3_axi_wlast   ),
    .s3_axi_wvalid  ( s3_axi_wvalid  ),
    .s3_axi_wready  ( s3_axi_wready  ),
    .s3_axi_bid     ( s3_axi_bid     ),
    .s3_axi_bresp   ( s3_axi_bresp   ),
    .s3_axi_bvalid  ( s3_axi_bvalid  ),
    .s3_axi_bready  ( s3_axi_bready  ),
    .m_awready      ( m_awready      ),
    .m_wready       ( m_wready       ),
    .m_bid          ( m_bid          ),
    .m_bresp        ( m_bresp        ),
    .m_bvalid       ( m_bvalid       ),
    .s_awid         ( s_awid         ),
    .s_awaddr       ( s_awaddr       ),
    .s_awlen        ( s_awlen        ),
    .s_awsize       ( s_awsize       ),
    .s_awburst      ( s_awburst      ),
    .s_awvalid      ( s_awvalid      ),
    .s_wdata        ( s_wdata        ),
    .s_wstrb        ( s_wstrb        ),
    .s_wlast        ( s_wlast        ),
    .s_wvalid       ( s_wvalid       ),
    .s_bready       ( s_bready       )
);
endmodule